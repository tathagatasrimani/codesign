
//------> /nfs/cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_wait_v1 (idat, rdy, ivld, dat, irdy, vld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  output             rdy;
  output             ivld;
  input  [width-1:0] dat;
  input              irdy;
  input              vld;

  wire   [width-1:0] idat;
  wire               rdy;
  wire               ivld;

  assign idat = dat;
  assign rdy = irdy;
  assign ivld = vld;

endmodule


//------> /nfs/cad/mentor/2019.11/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_out_wait_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_out_wait_v1 (dat, irdy, vld, idat, rdy, ivld);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] dat;
  output             irdy;
  output             vld;
  input  [width-1:0] idat;
  input              rdy;
  input              ivld;

  wire   [width-1:0] dat;
  wire               irdy;
  wire               vld;

  assign dat = idat;
  assign irdy = rdy;
  assign vld = ivld;

endmodule



//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   pmcewen@rsgvm14.stanford.edu
//  Generated date: Thu Feb 20 16:28:17 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    MatMult_run_run_fsm
//  FSM Module
// ------------------------------------------------------------------


module MatMult_run_run_fsm (
  clk, arst_n, run_wen, fsm_output, for_1_1_for_1_for_C_0_tr0
);
  input clk;
  input arst_n;
  input run_wen;
  output [3:0] fsm_output;
  reg [3:0] fsm_output;
  input for_1_1_for_1_for_C_0_tr0;


  // FSM State Type Declaration for MatMult_run_run_fsm_1
  parameter
    run_rlp_C_0 = 2'd0,
    main_C_0 = 2'd1,
    for_1_1_for_1_for_C_0 = 2'd2,
    main_C_1 = 2'd3;

  reg [1:0] state_var;
  reg [1:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : MatMult_run_run_fsm_1
    case (state_var)
      main_C_0 : begin
        fsm_output = 4'b0010;
        state_var_NS = for_1_1_for_1_for_C_0;
      end
      for_1_1_for_1_for_C_0 : begin
        fsm_output = 4'b0100;
        if ( for_1_1_for_1_for_C_0_tr0 ) begin
          state_var_NS = main_C_1;
        end
        else begin
          state_var_NS = for_1_1_for_1_for_C_0;
        end
      end
      main_C_1 : begin
        fsm_output = 4'b1000;
        state_var_NS = main_C_0;
      end
      // run_rlp_C_0
      default : begin
        fsm_output = 4'b0001;
        state_var_NS = main_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= run_rlp_C_0;
    end
    else if ( run_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_run_staller
// ------------------------------------------------------------------


module MatMult_run_staller (
  run_wen, a_chan_rsci_wen_comp, b_chan_rsci_wen_comp, c_chan_rsci_wen_comp
);
  output run_wen;
  input a_chan_rsci_wen_comp;
  input b_chan_rsci_wen_comp;
  input c_chan_rsci_wen_comp;



  // Interconnect Declarations for Component Instantiations 
  assign run_wen = a_chan_rsci_wen_comp & b_chan_rsci_wen_comp & c_chan_rsci_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_run_c_chan_rsci_c_chan_wait_dp
// ------------------------------------------------------------------


module MatMult_run_c_chan_rsci_c_chan_wait_dp (
  clk, arst_n, c_chan_rsci_oswt, c_chan_rsci_wen_comp, c_chan_rsci_biwt, c_chan_rsci_bdwt,
      c_chan_rsci_bcwt
);
  input clk;
  input arst_n;
  input c_chan_rsci_oswt;
  output c_chan_rsci_wen_comp;
  input c_chan_rsci_biwt;
  input c_chan_rsci_bdwt;
  output c_chan_rsci_bcwt;
  reg c_chan_rsci_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign c_chan_rsci_wen_comp = (~ c_chan_rsci_oswt) | c_chan_rsci_biwt | c_chan_rsci_bcwt;
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      c_chan_rsci_bcwt <= 1'b0;
    end
    else begin
      c_chan_rsci_bcwt <= ~((~(c_chan_rsci_bcwt | c_chan_rsci_biwt)) | c_chan_rsci_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_run_c_chan_rsci_c_chan_wait_ctrl
// ------------------------------------------------------------------


module MatMult_run_c_chan_rsci_c_chan_wait_ctrl (
  run_wen, c_chan_rsci_oswt, c_chan_rsci_irdy, c_chan_rsci_biwt, c_chan_rsci_bdwt,
      c_chan_rsci_bcwt, c_chan_rsci_ivld_run_sct
);
  input run_wen;
  input c_chan_rsci_oswt;
  input c_chan_rsci_irdy;
  output c_chan_rsci_biwt;
  output c_chan_rsci_bdwt;
  input c_chan_rsci_bcwt;
  output c_chan_rsci_ivld_run_sct;


  // Interconnect Declarations
  wire c_chan_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign c_chan_rsci_bdwt = c_chan_rsci_oswt & run_wen;
  assign c_chan_rsci_biwt = c_chan_rsci_ogwt & c_chan_rsci_irdy;
  assign c_chan_rsci_ogwt = c_chan_rsci_oswt & (~ c_chan_rsci_bcwt);
  assign c_chan_rsci_ivld_run_sct = c_chan_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_run_b_chan_rsci_b_chan_wait_dp
// ------------------------------------------------------------------


module MatMult_run_b_chan_rsci_b_chan_wait_dp (
  clk, arst_n, b_chan_rsci_oswt, b_chan_rsci_wen_comp, b_chan_rsci_idat_mxwt, b_chan_rsci_biwt,
      b_chan_rsci_bdwt, b_chan_rsci_bcwt, b_chan_rsci_idat
);
  input clk;
  input arst_n;
  input b_chan_rsci_oswt;
  output b_chan_rsci_wen_comp;
  output [399:0] b_chan_rsci_idat_mxwt;
  input b_chan_rsci_biwt;
  input b_chan_rsci_bdwt;
  output b_chan_rsci_bcwt;
  reg b_chan_rsci_bcwt;
  input [399:0] b_chan_rsci_idat;


  // Interconnect Declarations
  reg [399:0] b_chan_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign b_chan_rsci_wen_comp = (~ b_chan_rsci_oswt) | b_chan_rsci_biwt | b_chan_rsci_bcwt;
  assign b_chan_rsci_idat_mxwt = MUX_v_400_2_2(b_chan_rsci_idat, b_chan_rsci_idat_bfwt,
      b_chan_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      b_chan_rsci_bcwt <= 1'b0;
    end
    else begin
      b_chan_rsci_bcwt <= ~((~(b_chan_rsci_bcwt | b_chan_rsci_biwt)) | b_chan_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      b_chan_rsci_idat_bfwt <= 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ b_chan_rsci_bcwt ) begin
      b_chan_rsci_idat_bfwt <= b_chan_rsci_idat_mxwt;
    end
  end

  function automatic [399:0] MUX_v_400_2_2;
    input [399:0] input_0;
    input [399:0] input_1;
    input [0:0] sel;
    reg [399:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_400_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_run_b_chan_rsci_b_chan_wait_ctrl
// ------------------------------------------------------------------


module MatMult_run_b_chan_rsci_b_chan_wait_ctrl (
  run_wen, b_chan_rsci_oswt, b_chan_rsci_biwt, b_chan_rsci_bdwt, b_chan_rsci_bcwt,
      b_chan_rsci_irdy_run_sct, b_chan_rsci_ivld
);
  input run_wen;
  input b_chan_rsci_oswt;
  output b_chan_rsci_biwt;
  output b_chan_rsci_bdwt;
  input b_chan_rsci_bcwt;
  output b_chan_rsci_irdy_run_sct;
  input b_chan_rsci_ivld;


  // Interconnect Declarations
  wire b_chan_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign b_chan_rsci_bdwt = b_chan_rsci_oswt & run_wen;
  assign b_chan_rsci_biwt = b_chan_rsci_ogwt & b_chan_rsci_ivld;
  assign b_chan_rsci_ogwt = b_chan_rsci_oswt & (~ b_chan_rsci_bcwt);
  assign b_chan_rsci_irdy_run_sct = b_chan_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_run_a_chan_rsci_a_chan_wait_dp
// ------------------------------------------------------------------


module MatMult_run_a_chan_rsci_a_chan_wait_dp (
  clk, arst_n, a_chan_rsci_oswt, a_chan_rsci_wen_comp, a_chan_rsci_idat_mxwt, a_chan_rsci_biwt,
      a_chan_rsci_bdwt, a_chan_rsci_bcwt, a_chan_rsci_idat
);
  input clk;
  input arst_n;
  input a_chan_rsci_oswt;
  output a_chan_rsci_wen_comp;
  output [399:0] a_chan_rsci_idat_mxwt;
  input a_chan_rsci_biwt;
  input a_chan_rsci_bdwt;
  output a_chan_rsci_bcwt;
  reg a_chan_rsci_bcwt;
  input [399:0] a_chan_rsci_idat;


  // Interconnect Declarations
  reg [399:0] a_chan_rsci_idat_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign a_chan_rsci_wen_comp = (~ a_chan_rsci_oswt) | a_chan_rsci_biwt | a_chan_rsci_bcwt;
  assign a_chan_rsci_idat_mxwt = MUX_v_400_2_2(a_chan_rsci_idat, a_chan_rsci_idat_bfwt,
      a_chan_rsci_bcwt);
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      a_chan_rsci_bcwt <= 1'b0;
    end
    else begin
      a_chan_rsci_bcwt <= ~((~(a_chan_rsci_bcwt | a_chan_rsci_biwt)) | a_chan_rsci_bdwt);
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      a_chan_rsci_idat_bfwt <= 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ a_chan_rsci_bcwt ) begin
      a_chan_rsci_idat_bfwt <= a_chan_rsci_idat_mxwt;
    end
  end

  function automatic [399:0] MUX_v_400_2_2;
    input [399:0] input_0;
    input [399:0] input_1;
    input [0:0] sel;
    reg [399:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_400_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_run_a_chan_rsci_a_chan_wait_ctrl
// ------------------------------------------------------------------


module MatMult_run_a_chan_rsci_a_chan_wait_ctrl (
  run_wen, a_chan_rsci_oswt, a_chan_rsci_biwt, a_chan_rsci_bdwt, a_chan_rsci_bcwt,
      a_chan_rsci_irdy_run_sct, a_chan_rsci_ivld
);
  input run_wen;
  input a_chan_rsci_oswt;
  output a_chan_rsci_biwt;
  output a_chan_rsci_bdwt;
  input a_chan_rsci_bcwt;
  output a_chan_rsci_irdy_run_sct;
  input a_chan_rsci_ivld;


  // Interconnect Declarations
  wire a_chan_rsci_ogwt;


  // Interconnect Declarations for Component Instantiations 
  assign a_chan_rsci_bdwt = a_chan_rsci_oswt & run_wen;
  assign a_chan_rsci_biwt = a_chan_rsci_ogwt & a_chan_rsci_ivld;
  assign a_chan_rsci_ogwt = a_chan_rsci_oswt & (~ a_chan_rsci_bcwt);
  assign a_chan_rsci_irdy_run_sct = a_chan_rsci_ogwt;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_run_c_chan_rsci
// ------------------------------------------------------------------


module MatMult_run_c_chan_rsci (
  clk, arst_n, c_chan_rsc_dat, c_chan_rsc_vld, c_chan_rsc_rdy, run_wen, c_chan_rsci_oswt,
      c_chan_rsci_wen_comp, c_chan_rsci_idat
);
  input clk;
  input arst_n;
  output [399:0] c_chan_rsc_dat;
  output c_chan_rsc_vld;
  input c_chan_rsc_rdy;
  input run_wen;
  input c_chan_rsci_oswt;
  output c_chan_rsci_wen_comp;
  input [399:0] c_chan_rsci_idat;


  // Interconnect Declarations
  wire c_chan_rsci_irdy;
  wire c_chan_rsci_biwt;
  wire c_chan_rsci_bdwt;
  wire c_chan_rsci_bcwt;
  wire c_chan_rsci_ivld_run_sct;


  // Interconnect Declarations for Component Instantiations 
  ccs_out_wait_v1 #(.rscid(32'sd3),
  .width(32'sd400)) c_chan_rsci (
      .irdy(c_chan_rsci_irdy),
      .ivld(c_chan_rsci_ivld_run_sct),
      .idat(c_chan_rsci_idat),
      .rdy(c_chan_rsc_rdy),
      .vld(c_chan_rsc_vld),
      .dat(c_chan_rsc_dat)
    );
  MatMult_run_c_chan_rsci_c_chan_wait_ctrl MatMult_run_c_chan_rsci_c_chan_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .c_chan_rsci_oswt(c_chan_rsci_oswt),
      .c_chan_rsci_irdy(c_chan_rsci_irdy),
      .c_chan_rsci_biwt(c_chan_rsci_biwt),
      .c_chan_rsci_bdwt(c_chan_rsci_bdwt),
      .c_chan_rsci_bcwt(c_chan_rsci_bcwt),
      .c_chan_rsci_ivld_run_sct(c_chan_rsci_ivld_run_sct)
    );
  MatMult_run_c_chan_rsci_c_chan_wait_dp MatMult_run_c_chan_rsci_c_chan_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .c_chan_rsci_oswt(c_chan_rsci_oswt),
      .c_chan_rsci_wen_comp(c_chan_rsci_wen_comp),
      .c_chan_rsci_biwt(c_chan_rsci_biwt),
      .c_chan_rsci_bdwt(c_chan_rsci_bdwt),
      .c_chan_rsci_bcwt(c_chan_rsci_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_run_b_chan_rsci
// ------------------------------------------------------------------


module MatMult_run_b_chan_rsci (
  clk, arst_n, b_chan_rsc_dat, b_chan_rsc_vld, b_chan_rsc_rdy, run_wen, b_chan_rsci_oswt,
      b_chan_rsci_wen_comp, b_chan_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [399:0] b_chan_rsc_dat;
  input b_chan_rsc_vld;
  output b_chan_rsc_rdy;
  input run_wen;
  input b_chan_rsci_oswt;
  output b_chan_rsci_wen_comp;
  output [399:0] b_chan_rsci_idat_mxwt;


  // Interconnect Declarations
  wire b_chan_rsci_biwt;
  wire b_chan_rsci_bdwt;
  wire b_chan_rsci_bcwt;
  wire b_chan_rsci_irdy_run_sct;
  wire b_chan_rsci_ivld;
  wire [399:0] b_chan_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd2),
  .width(32'sd400)) b_chan_rsci (
      .rdy(b_chan_rsc_rdy),
      .vld(b_chan_rsc_vld),
      .dat(b_chan_rsc_dat),
      .irdy(b_chan_rsci_irdy_run_sct),
      .ivld(b_chan_rsci_ivld),
      .idat(b_chan_rsci_idat)
    );
  MatMult_run_b_chan_rsci_b_chan_wait_ctrl MatMult_run_b_chan_rsci_b_chan_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .b_chan_rsci_oswt(b_chan_rsci_oswt),
      .b_chan_rsci_biwt(b_chan_rsci_biwt),
      .b_chan_rsci_bdwt(b_chan_rsci_bdwt),
      .b_chan_rsci_bcwt(b_chan_rsci_bcwt),
      .b_chan_rsci_irdy_run_sct(b_chan_rsci_irdy_run_sct),
      .b_chan_rsci_ivld(b_chan_rsci_ivld)
    );
  MatMult_run_b_chan_rsci_b_chan_wait_dp MatMult_run_b_chan_rsci_b_chan_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .b_chan_rsci_oswt(b_chan_rsci_oswt),
      .b_chan_rsci_wen_comp(b_chan_rsci_wen_comp),
      .b_chan_rsci_idat_mxwt(b_chan_rsci_idat_mxwt),
      .b_chan_rsci_biwt(b_chan_rsci_biwt),
      .b_chan_rsci_bdwt(b_chan_rsci_bdwt),
      .b_chan_rsci_bcwt(b_chan_rsci_bcwt),
      .b_chan_rsci_idat(b_chan_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_run_a_chan_rsci
// ------------------------------------------------------------------


module MatMult_run_a_chan_rsci (
  clk, arst_n, a_chan_rsc_dat, a_chan_rsc_vld, a_chan_rsc_rdy, run_wen, a_chan_rsci_oswt,
      a_chan_rsci_wen_comp, a_chan_rsci_idat_mxwt
);
  input clk;
  input arst_n;
  input [399:0] a_chan_rsc_dat;
  input a_chan_rsc_vld;
  output a_chan_rsc_rdy;
  input run_wen;
  input a_chan_rsci_oswt;
  output a_chan_rsci_wen_comp;
  output [399:0] a_chan_rsci_idat_mxwt;


  // Interconnect Declarations
  wire a_chan_rsci_biwt;
  wire a_chan_rsci_bdwt;
  wire a_chan_rsci_bcwt;
  wire a_chan_rsci_irdy_run_sct;
  wire a_chan_rsci_ivld;
  wire [399:0] a_chan_rsci_idat;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_wait_v1 #(.rscid(32'sd1),
  .width(32'sd400)) a_chan_rsci (
      .rdy(a_chan_rsc_rdy),
      .vld(a_chan_rsc_vld),
      .dat(a_chan_rsc_dat),
      .irdy(a_chan_rsci_irdy_run_sct),
      .ivld(a_chan_rsci_ivld),
      .idat(a_chan_rsci_idat)
    );
  MatMult_run_a_chan_rsci_a_chan_wait_ctrl MatMult_run_a_chan_rsci_a_chan_wait_ctrl_inst
      (
      .run_wen(run_wen),
      .a_chan_rsci_oswt(a_chan_rsci_oswt),
      .a_chan_rsci_biwt(a_chan_rsci_biwt),
      .a_chan_rsci_bdwt(a_chan_rsci_bdwt),
      .a_chan_rsci_bcwt(a_chan_rsci_bcwt),
      .a_chan_rsci_irdy_run_sct(a_chan_rsci_irdy_run_sct),
      .a_chan_rsci_ivld(a_chan_rsci_ivld)
    );
  MatMult_run_a_chan_rsci_a_chan_wait_dp MatMult_run_a_chan_rsci_a_chan_wait_dp_inst
      (
      .clk(clk),
      .arst_n(arst_n),
      .a_chan_rsci_oswt(a_chan_rsci_oswt),
      .a_chan_rsci_wen_comp(a_chan_rsci_wen_comp),
      .a_chan_rsci_idat_mxwt(a_chan_rsci_idat_mxwt),
      .a_chan_rsci_biwt(a_chan_rsci_biwt),
      .a_chan_rsci_bdwt(a_chan_rsci_bdwt),
      .a_chan_rsci_bcwt(a_chan_rsci_bcwt),
      .a_chan_rsci_idat(a_chan_rsci_idat)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_run
// ------------------------------------------------------------------


module MatMult_run (
  clk, arst_n, a_chan_rsc_dat, a_chan_rsc_vld, a_chan_rsc_rdy, b_chan_rsc_dat, b_chan_rsc_vld,
      b_chan_rsc_rdy, c_chan_rsc_dat, c_chan_rsc_vld, c_chan_rsc_rdy
);
  input clk;
  input arst_n;
  input [399:0] a_chan_rsc_dat;
  input a_chan_rsc_vld;
  output a_chan_rsc_rdy;
  input [399:0] b_chan_rsc_dat;
  input b_chan_rsc_vld;
  output b_chan_rsc_rdy;
  output [399:0] c_chan_rsc_dat;
  output c_chan_rsc_vld;
  input c_chan_rsc_rdy;


  // Interconnect Declarations
  wire run_wen;
  wire a_chan_rsci_wen_comp;
  wire [399:0] a_chan_rsci_idat_mxwt;
  wire b_chan_rsci_wen_comp;
  wire [399:0] b_chan_rsci_idat_mxwt;
  wire c_chan_rsci_wen_comp;
  reg [15:0] c_chan_rsci_idat_399_384;
  reg [15:0] c_chan_rsci_idat_383_368;
  reg [15:0] c_chan_rsci_idat_367_352;
  reg [15:0] c_chan_rsci_idat_351_336;
  reg [15:0] c_chan_rsci_idat_335_320;
  reg [15:0] c_chan_rsci_idat_319_304;
  reg [15:0] c_chan_rsci_idat_303_288;
  reg [15:0] c_chan_rsci_idat_287_272;
  reg [15:0] c_chan_rsci_idat_271_256;
  reg [15:0] c_chan_rsci_idat_255_240;
  reg [15:0] c_chan_rsci_idat_239_224;
  reg [15:0] c_chan_rsci_idat_223_208;
  reg [15:0] c_chan_rsci_idat_207_192;
  reg [15:0] c_chan_rsci_idat_191_176;
  reg [15:0] c_chan_rsci_idat_175_160;
  reg [15:0] c_chan_rsci_idat_159_144;
  reg [15:0] c_chan_rsci_idat_143_128;
  reg [15:0] c_chan_rsci_idat_127_112;
  reg [15:0] c_chan_rsci_idat_111_96;
  reg [15:0] c_chan_rsci_idat_95_80;
  reg [15:0] c_chan_rsci_idat_79_64;
  reg [15:0] c_chan_rsci_idat_63_48;
  reg [15:0] c_chan_rsci_idat_47_32;
  reg [15:0] c_chan_rsci_idat_31_16;
  reg [15:0] c_chan_rsci_idat_15_0;
  wire [3:0] fsm_output;
  wire for_1_for_for_and_21_tmp;
  wire c_chan_and_cse;
  reg reg_c_chan_rsci_ivld_run_psct_cse;
  reg reg_b_chan_rsci_irdy_run_psct_cse;
  reg [399:0] a_value_value_sva;
  reg [399:0] b_value_value_sva;
  reg [15:0] for_1_for_tmp_9_sva;
  reg [2:0] for_1_for_for_k_2_0_9_sva;
  reg [15:0] for_1_for_tmp_13_sva;
  reg [2:0] for_1_for_for_k_2_0_13_sva;
  reg [15:0] for_1_for_tmp_17_sva;
  reg [2:0] for_1_for_for_k_2_0_17_sva;
  reg [15:0] for_1_for_tmp_21_sva;
  reg [2:0] for_1_for_for_k_2_0_21_sva;
  reg [15:0] for_1_for_tmp_5_sva;
  reg [2:0] for_1_for_for_k_2_0_5_sva;
  reg [15:0] for_1_for_tmp_10_sva;
  reg [2:0] for_1_for_for_k_2_0_10_sva;
  reg [15:0] for_1_for_tmp_14_sva;
  reg [2:0] for_1_for_for_k_2_0_14_sva;
  reg [15:0] for_1_for_tmp_18_sva;
  reg [2:0] for_1_for_for_k_2_0_18_sva;
  reg [15:0] for_1_for_tmp_22_sva;
  reg [2:0] for_1_for_for_k_2_0_22_sva;
  reg [15:0] for_1_for_tmp_6_sva;
  reg [2:0] for_1_for_for_k_2_0_6_sva;
  reg [15:0] for_1_for_tmp_11_sva;
  reg [2:0] for_1_for_for_k_2_0_11_sva;
  reg [15:0] for_1_for_tmp_15_sva;
  reg [2:0] for_1_for_for_k_2_0_15_sva;
  reg [15:0] for_1_for_tmp_19_sva;
  reg [2:0] for_1_for_for_k_2_0_19_sva;
  reg [15:0] for_1_for_tmp_23_sva;
  reg [2:0] for_1_for_for_k_2_0_23_sva;
  reg [15:0] for_1_for_tmp_7_sva;
  reg [2:0] for_1_for_for_k_2_0_7_sva;
  reg [15:0] for_1_for_tmp_12_sva;
  reg [2:0] for_1_for_for_k_2_0_12_sva;
  reg [15:0] for_1_for_tmp_16_sva;
  reg [2:0] for_1_for_for_k_2_0_16_sva;
  reg [15:0] for_1_for_tmp_20_sva;
  reg [2:0] for_1_for_for_k_2_0_20_sva;
  reg [15:0] for_1_for_tmp_24_sva;
  reg [2:0] for_1_for_for_k_2_0_24_sva;
  reg [15:0] for_1_for_tmp_8_sva;
  reg [2:0] for_1_for_for_k_2_0_8_sva;
  reg [15:0] for_1_for_tmp_1_sva;
  reg [2:0] for_1_for_for_k_2_0_1_sva;
  reg [15:0] for_1_for_tmp_2_sva;
  reg [2:0] for_1_for_for_k_2_0_2_sva;
  reg [15:0] for_1_for_tmp_3_sva;
  reg [2:0] for_1_for_for_k_2_0_3_sva;
  reg [15:0] for_1_for_tmp_4_sva;
  reg [2:0] for_1_for_for_k_2_0_4_sva;
  reg [15:0] for_1_for_tmp_sva;
  reg [2:0] for_1_for_for_k_2_0_sva;
  wire [15:0] for_1_for_tmp_9_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_9_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_13_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_13_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_17_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_17_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_21_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_21_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_5_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_5_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_10_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_10_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_14_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_14_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_18_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_18_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_22_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_22_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_6_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_6_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_11_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_11_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_15_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_15_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_19_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_19_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_23_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_23_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_7_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_7_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_12_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_12_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_16_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_16_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_20_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_20_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_24_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_24_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_8_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_8_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_1_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_1_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_2_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_2_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_3_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_3_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_4_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_4_sva_1_mx0w0;
  wire [15:0] for_1_for_tmp_sva_1_mx0w0;
  wire [16:0] nl_for_1_for_tmp_sva_1_mx0w0;
  wire [2:0] for_1_for_for_k_2_0_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_sva_2;
  wire [2:0] for_1_for_for_k_2_0_4_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_4_sva_2;
  wire [2:0] for_1_for_for_k_2_0_3_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_3_sva_2;
  wire [2:0] for_1_for_for_k_2_0_2_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_2_sva_2;
  wire [2:0] for_1_for_for_k_2_0_1_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_1_sva_2;
  wire [2:0] for_1_for_for_k_2_0_8_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_8_sva_2;
  wire [2:0] for_1_for_for_k_2_0_24_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_24_sva_2;
  wire [2:0] for_1_for_for_k_2_0_20_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_20_sva_2;
  wire [2:0] for_1_for_for_k_2_0_16_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_16_sva_2;
  wire [2:0] for_1_for_for_k_2_0_12_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_12_sva_2;
  wire [2:0] for_1_for_for_k_2_0_7_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_7_sva_2;
  wire [2:0] for_1_for_for_k_2_0_23_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_23_sva_2;
  wire [2:0] for_1_for_for_k_2_0_19_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_19_sva_2;
  wire [2:0] for_1_for_for_k_2_0_15_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_15_sva_2;
  wire [2:0] for_1_for_for_k_2_0_11_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_11_sva_2;
  wire [2:0] for_1_for_for_k_2_0_6_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_6_sva_2;
  wire [2:0] for_1_for_for_k_2_0_22_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_22_sva_2;
  wire [2:0] for_1_for_for_k_2_0_18_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_18_sva_2;
  wire [2:0] for_1_for_for_k_2_0_14_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_14_sva_2;
  wire [2:0] for_1_for_for_k_2_0_10_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_10_sva_2;
  wire [2:0] for_1_for_for_k_2_0_5_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_5_sva_2;
  wire [2:0] for_1_for_for_k_2_0_21_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_21_sva_2;
  wire [2:0] for_1_for_for_k_2_0_17_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_17_sva_2;
  wire [2:0] for_1_for_for_k_2_0_13_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_13_sva_2;
  wire [2:0] for_1_for_for_k_2_0_9_sva_2;
  wire [3:0] nl_for_1_for_for_k_2_0_9_sva_2;
  wire [15:0] for_1_5_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1;
  wire [15:0] for_1_1_for_5_for_slc_b_value_value_16_15_0_ncse_sva_1;
  wire [15:0] for_1_1_for_4_for_slc_b_value_value_16_15_0_ncse_sva_1;
  wire [15:0] for_1_1_for_3_for_slc_b_value_value_16_15_0_ncse_sva_1;
  wire [15:0] for_1_1_for_2_for_slc_b_value_value_16_15_0_ncse_sva_1;
  wire [15:0] for_1_1_for_1_for_slc_b_value_value_16_15_0_ncse_sva_1;
  wire [15:0] for_1_4_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1;
  wire [15:0] for_1_3_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1;
  wire [15:0] for_1_2_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1;
  wire [15:0] for_1_1_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1;
  wire [2:0] for_1_for_for_acc_18_psp_1;
  wire [3:0] nl_for_1_for_for_acc_18_psp_1;
  wire a_value_value_and_cse;

  wire[15:0] for_1_1_for_1_for_mul_nl;
  wire signed [31:0] nl_for_1_1_for_1_for_mul_nl;
  wire[15:0] for_1_1_for_2_for_mul_nl;
  wire signed [31:0] nl_for_1_1_for_2_for_mul_nl;
  wire[15:0] for_1_1_for_3_for_mul_nl;
  wire signed [31:0] nl_for_1_1_for_3_for_mul_nl;
  wire[15:0] for_1_1_for_4_for_mul_nl;
  wire signed [31:0] nl_for_1_1_for_4_for_mul_nl;
  wire[15:0] for_1_1_for_5_for_mul_nl;
  wire signed [31:0] nl_for_1_1_for_5_for_mul_nl;
  wire[15:0] for_1_2_for_1_for_mul_nl;
  wire signed [31:0] nl_for_1_2_for_1_for_mul_nl;
  wire[15:0] for_1_2_for_2_for_mul_nl;
  wire signed [31:0] nl_for_1_2_for_2_for_mul_nl;
  wire[15:0] for_1_2_for_3_for_mul_nl;
  wire signed [31:0] nl_for_1_2_for_3_for_mul_nl;
  wire[15:0] for_1_2_for_4_for_mul_nl;
  wire signed [31:0] nl_for_1_2_for_4_for_mul_nl;
  wire[15:0] for_1_2_for_5_for_mul_nl;
  wire signed [31:0] nl_for_1_2_for_5_for_mul_nl;
  wire[15:0] for_1_3_for_1_for_mul_nl;
  wire signed [31:0] nl_for_1_3_for_1_for_mul_nl;
  wire[15:0] for_1_3_for_2_for_mul_nl;
  wire signed [31:0] nl_for_1_3_for_2_for_mul_nl;
  wire[15:0] for_1_3_for_3_for_mul_nl;
  wire signed [31:0] nl_for_1_3_for_3_for_mul_nl;
  wire[15:0] for_1_3_for_4_for_mul_nl;
  wire signed [31:0] nl_for_1_3_for_4_for_mul_nl;
  wire[15:0] for_1_3_for_5_for_mul_nl;
  wire signed [31:0] nl_for_1_3_for_5_for_mul_nl;
  wire[15:0] for_1_4_for_1_for_mul_nl;
  wire signed [31:0] nl_for_1_4_for_1_for_mul_nl;
  wire[15:0] for_1_4_for_2_for_mul_nl;
  wire signed [31:0] nl_for_1_4_for_2_for_mul_nl;
  wire[15:0] for_1_4_for_3_for_mul_nl;
  wire signed [31:0] nl_for_1_4_for_3_for_mul_nl;
  wire[15:0] for_1_4_for_4_for_mul_nl;
  wire signed [31:0] nl_for_1_4_for_4_for_mul_nl;
  wire[15:0] for_1_4_for_5_for_mul_nl;
  wire signed [31:0] nl_for_1_4_for_5_for_mul_nl;
  wire[15:0] for_1_5_for_1_for_mul_nl;
  wire signed [31:0] nl_for_1_5_for_1_for_mul_nl;
  wire[15:0] for_1_5_for_2_for_mul_nl;
  wire signed [31:0] nl_for_1_5_for_2_for_mul_nl;
  wire[15:0] for_1_5_for_3_for_mul_nl;
  wire signed [31:0] nl_for_1_5_for_3_for_mul_nl;
  wire[15:0] for_1_5_for_4_for_mul_nl;
  wire signed [31:0] nl_for_1_5_for_4_for_mul_nl;
  wire[15:0] for_1_5_for_5_for_mul_nl;
  wire signed [31:0] nl_for_1_5_for_5_for_mul_nl;
  wire[2:0] for_1_1_for_for_acc_7_nl;
  wire[4:0] nl_for_1_1_for_for_acc_7_nl;
  wire[2:0] for_1_for_for_acc_19_nl;
  wire[3:0] nl_for_1_for_for_acc_19_nl;
  wire[3:0] for_1_1_for_for_acc_nl;
  wire[5:0] nl_for_1_1_for_for_acc_nl;
  wire[4:0] for_1_1_for_2_for_acc_6_nl;
  wire[6:0] nl_for_1_1_for_2_for_acc_6_nl;
  wire[2:0] for_1_1_for_for_acc_8_nl;
  wire[3:0] nl_for_1_1_for_for_acc_8_nl;
  wire[2:0] for_1_4_for_1_for_acc_5_nl;
  wire[3:0] nl_for_1_4_for_1_for_acc_5_nl;
  wire[1:0] for_1_for_for_acc_nl;
  wire[2:0] nl_for_1_for_for_acc_nl;
  wire[2:0] for_1_2_for_1_for_acc_5_nl;
  wire[3:0] nl_for_1_2_for_1_for_acc_5_nl;
  wire[3:0] for_1_1_for_1_for_acc_nl;
  wire[4:0] nl_for_1_1_for_1_for_acc_nl;
  wire[3:0] for_1_1_for_2_for_acc_nl;
  wire[4:0] nl_for_1_1_for_2_for_acc_nl;
  wire[3:0] for_1_1_for_3_for_acc_nl;
  wire[4:0] nl_for_1_1_for_3_for_acc_nl;
  wire[3:0] for_1_1_for_4_for_acc_nl;
  wire[4:0] nl_for_1_1_for_4_for_acc_nl;
  wire[3:0] for_1_1_for_5_for_acc_nl;
  wire[4:0] nl_for_1_1_for_5_for_acc_nl;
  wire[3:0] for_1_2_for_1_for_acc_nl;
  wire[4:0] nl_for_1_2_for_1_for_acc_nl;
  wire[3:0] for_1_2_for_2_for_acc_nl;
  wire[4:0] nl_for_1_2_for_2_for_acc_nl;
  wire[3:0] for_1_2_for_3_for_acc_nl;
  wire[4:0] nl_for_1_2_for_3_for_acc_nl;
  wire[3:0] for_1_2_for_4_for_acc_nl;
  wire[4:0] nl_for_1_2_for_4_for_acc_nl;
  wire[3:0] for_1_2_for_5_for_acc_nl;
  wire[4:0] nl_for_1_2_for_5_for_acc_nl;
  wire[3:0] for_1_3_for_1_for_acc_nl;
  wire[4:0] nl_for_1_3_for_1_for_acc_nl;
  wire[3:0] for_1_3_for_2_for_acc_nl;
  wire[4:0] nl_for_1_3_for_2_for_acc_nl;
  wire[3:0] for_1_3_for_3_for_acc_nl;
  wire[4:0] nl_for_1_3_for_3_for_acc_nl;
  wire[3:0] for_1_3_for_4_for_acc_nl;
  wire[4:0] nl_for_1_3_for_4_for_acc_nl;
  wire[3:0] for_1_3_for_5_for_acc_nl;
  wire[4:0] nl_for_1_3_for_5_for_acc_nl;
  wire[3:0] for_1_4_for_1_for_acc_nl;
  wire[4:0] nl_for_1_4_for_1_for_acc_nl;
  wire[3:0] for_1_4_for_2_for_acc_nl;
  wire[4:0] nl_for_1_4_for_2_for_acc_nl;
  wire[3:0] for_1_4_for_3_for_acc_nl;
  wire[4:0] nl_for_1_4_for_3_for_acc_nl;
  wire[3:0] for_1_4_for_4_for_acc_nl;
  wire[4:0] nl_for_1_4_for_4_for_acc_nl;
  wire[3:0] for_1_4_for_5_for_acc_nl;
  wire[4:0] nl_for_1_4_for_5_for_acc_nl;
  wire[3:0] for_1_5_for_1_for_acc_nl;
  wire[4:0] nl_for_1_5_for_1_for_acc_nl;
  wire[3:0] for_1_5_for_2_for_acc_nl;
  wire[4:0] nl_for_1_5_for_2_for_acc_nl;
  wire[3:0] for_1_5_for_3_for_acc_nl;
  wire[4:0] nl_for_1_5_for_3_for_acc_nl;
  wire[3:0] for_1_5_for_4_for_acc_nl;
  wire[4:0] nl_for_1_5_for_4_for_acc_nl;
  wire[3:0] for_1_5_for_5_for_acc_nl;
  wire[4:0] nl_for_1_5_for_5_for_acc_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [399:0] nl_MatMult_run_c_chan_rsci_inst_c_chan_rsci_idat;
  assign nl_MatMult_run_c_chan_rsci_inst_c_chan_rsci_idat = {c_chan_rsci_idat_399_384
      , c_chan_rsci_idat_383_368 , c_chan_rsci_idat_367_352 , c_chan_rsci_idat_351_336
      , c_chan_rsci_idat_335_320 , c_chan_rsci_idat_319_304 , c_chan_rsci_idat_303_288
      , c_chan_rsci_idat_287_272 , c_chan_rsci_idat_271_256 , c_chan_rsci_idat_255_240
      , c_chan_rsci_idat_239_224 , c_chan_rsci_idat_223_208 , c_chan_rsci_idat_207_192
      , c_chan_rsci_idat_191_176 , c_chan_rsci_idat_175_160 , c_chan_rsci_idat_159_144
      , c_chan_rsci_idat_143_128 , c_chan_rsci_idat_127_112 , c_chan_rsci_idat_111_96
      , c_chan_rsci_idat_95_80 , c_chan_rsci_idat_79_64 , c_chan_rsci_idat_63_48
      , c_chan_rsci_idat_47_32 , c_chan_rsci_idat_31_16 , c_chan_rsci_idat_15_0};
  MatMult_run_a_chan_rsci MatMult_run_a_chan_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .a_chan_rsc_dat(a_chan_rsc_dat),
      .a_chan_rsc_vld(a_chan_rsc_vld),
      .a_chan_rsc_rdy(a_chan_rsc_rdy),
      .run_wen(run_wen),
      .a_chan_rsci_oswt(reg_b_chan_rsci_irdy_run_psct_cse),
      .a_chan_rsci_wen_comp(a_chan_rsci_wen_comp),
      .a_chan_rsci_idat_mxwt(a_chan_rsci_idat_mxwt)
    );
  MatMult_run_b_chan_rsci MatMult_run_b_chan_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .b_chan_rsc_dat(b_chan_rsc_dat),
      .b_chan_rsc_vld(b_chan_rsc_vld),
      .b_chan_rsc_rdy(b_chan_rsc_rdy),
      .run_wen(run_wen),
      .b_chan_rsci_oswt(reg_b_chan_rsci_irdy_run_psct_cse),
      .b_chan_rsci_wen_comp(b_chan_rsci_wen_comp),
      .b_chan_rsci_idat_mxwt(b_chan_rsci_idat_mxwt)
    );
  MatMult_run_c_chan_rsci MatMult_run_c_chan_rsci_inst (
      .clk(clk),
      .arst_n(arst_n),
      .c_chan_rsc_dat(c_chan_rsc_dat),
      .c_chan_rsc_vld(c_chan_rsc_vld),
      .c_chan_rsc_rdy(c_chan_rsc_rdy),
      .run_wen(run_wen),
      .c_chan_rsci_oswt(reg_c_chan_rsci_ivld_run_psct_cse),
      .c_chan_rsci_wen_comp(c_chan_rsci_wen_comp),
      .c_chan_rsci_idat(nl_MatMult_run_c_chan_rsci_inst_c_chan_rsci_idat[399:0])
    );
  MatMult_run_staller MatMult_run_staller_inst (
      .run_wen(run_wen),
      .a_chan_rsci_wen_comp(a_chan_rsci_wen_comp),
      .b_chan_rsci_wen_comp(b_chan_rsci_wen_comp),
      .c_chan_rsci_wen_comp(c_chan_rsci_wen_comp)
    );
  MatMult_run_run_fsm MatMult_run_run_fsm_inst (
      .clk(clk),
      .arst_n(arst_n),
      .run_wen(run_wen),
      .fsm_output(fsm_output),
      .for_1_1_for_1_for_C_0_tr0(for_1_for_for_and_21_tmp)
    );
  assign c_chan_and_cse = run_wen & (fsm_output[2]) & for_1_for_for_and_21_tmp;
  assign a_value_value_and_cse = run_wen & (~ (fsm_output[2]));
  assign nl_for_1_1_for_1_for_mul_nl = $signed(for_1_1_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_1_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_1_for_1_for_mul_nl = nl_for_1_1_for_1_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_9_sva_1_mx0w0 = for_1_for_tmp_9_sva + (for_1_1_for_1_for_mul_nl);
  assign for_1_for_tmp_9_sva_1_mx0w0 = nl_for_1_for_tmp_9_sva_1_mx0w0[15:0];
  assign nl_for_1_1_for_2_for_mul_nl = $signed(for_1_1_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_2_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_1_for_2_for_mul_nl = nl_for_1_1_for_2_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_13_sva_1_mx0w0 = for_1_for_tmp_13_sva + (for_1_1_for_2_for_mul_nl);
  assign for_1_for_tmp_13_sva_1_mx0w0 = nl_for_1_for_tmp_13_sva_1_mx0w0[15:0];
  assign nl_for_1_1_for_3_for_mul_nl = $signed(for_1_1_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_3_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_1_for_3_for_mul_nl = nl_for_1_1_for_3_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_17_sva_1_mx0w0 = for_1_for_tmp_17_sva + (for_1_1_for_3_for_mul_nl);
  assign for_1_for_tmp_17_sva_1_mx0w0 = nl_for_1_for_tmp_17_sva_1_mx0w0[15:0];
  assign nl_for_1_1_for_4_for_mul_nl = $signed(for_1_1_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_4_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_1_for_4_for_mul_nl = nl_for_1_1_for_4_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_21_sva_1_mx0w0 = for_1_for_tmp_21_sva + (for_1_1_for_4_for_mul_nl);
  assign for_1_for_tmp_21_sva_1_mx0w0 = nl_for_1_for_tmp_21_sva_1_mx0w0[15:0];
  assign nl_for_1_1_for_5_for_mul_nl = $signed(for_1_1_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_5_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_1_for_5_for_mul_nl = nl_for_1_1_for_5_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_5_sva_1_mx0w0 = for_1_for_tmp_5_sva + (for_1_1_for_5_for_mul_nl);
  assign for_1_for_tmp_5_sva_1_mx0w0 = nl_for_1_for_tmp_5_sva_1_mx0w0[15:0];
  assign nl_for_1_2_for_1_for_mul_nl = $signed(for_1_2_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_1_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_2_for_1_for_mul_nl = nl_for_1_2_for_1_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_10_sva_1_mx0w0 = for_1_for_tmp_10_sva + (for_1_2_for_1_for_mul_nl);
  assign for_1_for_tmp_10_sva_1_mx0w0 = nl_for_1_for_tmp_10_sva_1_mx0w0[15:0];
  assign nl_for_1_2_for_2_for_mul_nl = $signed(for_1_2_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_2_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_2_for_2_for_mul_nl = nl_for_1_2_for_2_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_14_sva_1_mx0w0 = for_1_for_tmp_14_sva + (for_1_2_for_2_for_mul_nl);
  assign for_1_for_tmp_14_sva_1_mx0w0 = nl_for_1_for_tmp_14_sva_1_mx0w0[15:0];
  assign nl_for_1_2_for_3_for_mul_nl = $signed(for_1_2_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_3_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_2_for_3_for_mul_nl = nl_for_1_2_for_3_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_18_sva_1_mx0w0 = for_1_for_tmp_18_sva + (for_1_2_for_3_for_mul_nl);
  assign for_1_for_tmp_18_sva_1_mx0w0 = nl_for_1_for_tmp_18_sva_1_mx0w0[15:0];
  assign nl_for_1_2_for_4_for_mul_nl = $signed(for_1_2_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_4_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_2_for_4_for_mul_nl = nl_for_1_2_for_4_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_22_sva_1_mx0w0 = for_1_for_tmp_22_sva + (for_1_2_for_4_for_mul_nl);
  assign for_1_for_tmp_22_sva_1_mx0w0 = nl_for_1_for_tmp_22_sva_1_mx0w0[15:0];
  assign nl_for_1_2_for_5_for_mul_nl = $signed(for_1_2_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_5_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_2_for_5_for_mul_nl = nl_for_1_2_for_5_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_6_sva_1_mx0w0 = for_1_for_tmp_6_sva + (for_1_2_for_5_for_mul_nl);
  assign for_1_for_tmp_6_sva_1_mx0w0 = nl_for_1_for_tmp_6_sva_1_mx0w0[15:0];
  assign nl_for_1_3_for_1_for_mul_nl = $signed(for_1_3_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_1_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_3_for_1_for_mul_nl = nl_for_1_3_for_1_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_11_sva_1_mx0w0 = for_1_for_tmp_11_sva + (for_1_3_for_1_for_mul_nl);
  assign for_1_for_tmp_11_sva_1_mx0w0 = nl_for_1_for_tmp_11_sva_1_mx0w0[15:0];
  assign nl_for_1_3_for_2_for_mul_nl = $signed(for_1_3_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_2_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_3_for_2_for_mul_nl = nl_for_1_3_for_2_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_15_sva_1_mx0w0 = for_1_for_tmp_15_sva + (for_1_3_for_2_for_mul_nl);
  assign for_1_for_tmp_15_sva_1_mx0w0 = nl_for_1_for_tmp_15_sva_1_mx0w0[15:0];
  assign nl_for_1_3_for_3_for_mul_nl = $signed(for_1_3_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_3_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_3_for_3_for_mul_nl = nl_for_1_3_for_3_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_19_sva_1_mx0w0 = for_1_for_tmp_19_sva + (for_1_3_for_3_for_mul_nl);
  assign for_1_for_tmp_19_sva_1_mx0w0 = nl_for_1_for_tmp_19_sva_1_mx0w0[15:0];
  assign nl_for_1_3_for_4_for_mul_nl = $signed(for_1_3_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_4_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_3_for_4_for_mul_nl = nl_for_1_3_for_4_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_23_sva_1_mx0w0 = for_1_for_tmp_23_sva + (for_1_3_for_4_for_mul_nl);
  assign for_1_for_tmp_23_sva_1_mx0w0 = nl_for_1_for_tmp_23_sva_1_mx0w0[15:0];
  assign nl_for_1_3_for_5_for_mul_nl = $signed(for_1_3_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_5_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_3_for_5_for_mul_nl = nl_for_1_3_for_5_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_7_sva_1_mx0w0 = for_1_for_tmp_7_sva + (for_1_3_for_5_for_mul_nl);
  assign for_1_for_tmp_7_sva_1_mx0w0 = nl_for_1_for_tmp_7_sva_1_mx0w0[15:0];
  assign nl_for_1_4_for_1_for_mul_nl = $signed(for_1_4_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_1_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_4_for_1_for_mul_nl = nl_for_1_4_for_1_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_12_sva_1_mx0w0 = for_1_for_tmp_12_sva + (for_1_4_for_1_for_mul_nl);
  assign for_1_for_tmp_12_sva_1_mx0w0 = nl_for_1_for_tmp_12_sva_1_mx0w0[15:0];
  assign nl_for_1_4_for_2_for_mul_nl = $signed(for_1_4_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_2_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_4_for_2_for_mul_nl = nl_for_1_4_for_2_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_16_sva_1_mx0w0 = for_1_for_tmp_16_sva + (for_1_4_for_2_for_mul_nl);
  assign for_1_for_tmp_16_sva_1_mx0w0 = nl_for_1_for_tmp_16_sva_1_mx0w0[15:0];
  assign nl_for_1_4_for_3_for_mul_nl = $signed(for_1_4_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_3_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_4_for_3_for_mul_nl = nl_for_1_4_for_3_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_20_sva_1_mx0w0 = for_1_for_tmp_20_sva + (for_1_4_for_3_for_mul_nl);
  assign for_1_for_tmp_20_sva_1_mx0w0 = nl_for_1_for_tmp_20_sva_1_mx0w0[15:0];
  assign nl_for_1_4_for_4_for_mul_nl = $signed(for_1_4_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_4_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_4_for_4_for_mul_nl = nl_for_1_4_for_4_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_24_sva_1_mx0w0 = for_1_for_tmp_24_sva + (for_1_4_for_4_for_mul_nl);
  assign for_1_for_tmp_24_sva_1_mx0w0 = nl_for_1_for_tmp_24_sva_1_mx0w0[15:0];
  assign nl_for_1_4_for_5_for_mul_nl = $signed(for_1_4_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_5_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_4_for_5_for_mul_nl = nl_for_1_4_for_5_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_8_sva_1_mx0w0 = for_1_for_tmp_8_sva + (for_1_4_for_5_for_mul_nl);
  assign for_1_for_tmp_8_sva_1_mx0w0 = nl_for_1_for_tmp_8_sva_1_mx0w0[15:0];
  assign nl_for_1_5_for_1_for_mul_nl = $signed(for_1_5_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_1_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_5_for_1_for_mul_nl = nl_for_1_5_for_1_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_1_sva_1_mx0w0 = for_1_for_tmp_1_sva + (for_1_5_for_1_for_mul_nl);
  assign for_1_for_tmp_1_sva_1_mx0w0 = nl_for_1_for_tmp_1_sva_1_mx0w0[15:0];
  assign nl_for_1_5_for_2_for_mul_nl = $signed(for_1_5_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_2_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_5_for_2_for_mul_nl = nl_for_1_5_for_2_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_2_sva_1_mx0w0 = for_1_for_tmp_2_sva + (for_1_5_for_2_for_mul_nl);
  assign for_1_for_tmp_2_sva_1_mx0w0 = nl_for_1_for_tmp_2_sva_1_mx0w0[15:0];
  assign nl_for_1_5_for_3_for_mul_nl = $signed(for_1_5_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_3_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_5_for_3_for_mul_nl = nl_for_1_5_for_3_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_3_sva_1_mx0w0 = for_1_for_tmp_3_sva + (for_1_5_for_3_for_mul_nl);
  assign for_1_for_tmp_3_sva_1_mx0w0 = nl_for_1_for_tmp_3_sva_1_mx0w0[15:0];
  assign nl_for_1_5_for_4_for_mul_nl = $signed(for_1_5_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_4_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_5_for_4_for_mul_nl = nl_for_1_5_for_4_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_4_sva_1_mx0w0 = for_1_for_tmp_4_sva + (for_1_5_for_4_for_mul_nl);
  assign for_1_for_tmp_4_sva_1_mx0w0 = nl_for_1_for_tmp_4_sva_1_mx0w0[15:0];
  assign nl_for_1_5_for_5_for_mul_nl = $signed(for_1_5_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1)
      * $signed(for_1_1_for_5_for_slc_b_value_value_16_15_0_ncse_sva_1);
  assign for_1_5_for_5_for_mul_nl = nl_for_1_5_for_5_for_mul_nl[15:0];
  assign nl_for_1_for_tmp_sva_1_mx0w0 = for_1_for_tmp_sva + (for_1_5_for_5_for_mul_nl);
  assign for_1_for_tmp_sva_1_mx0w0 = nl_for_1_for_tmp_sva_1_mx0w0[15:0];
  assign nl_for_1_for_for_k_2_0_sva_2 = for_1_for_for_k_2_0_sva + 3'b001;
  assign for_1_for_for_k_2_0_sva_2 = nl_for_1_for_for_k_2_0_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_4_sva_2 = for_1_for_for_k_2_0_4_sva + 3'b001;
  assign for_1_for_for_k_2_0_4_sva_2 = nl_for_1_for_for_k_2_0_4_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_3_sva_2 = for_1_for_for_k_2_0_3_sva + 3'b001;
  assign for_1_for_for_k_2_0_3_sva_2 = nl_for_1_for_for_k_2_0_3_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_2_sva_2 = for_1_for_for_k_2_0_2_sva + 3'b001;
  assign for_1_for_for_k_2_0_2_sva_2 = nl_for_1_for_for_k_2_0_2_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_1_sva_2 = for_1_for_for_k_2_0_1_sva + 3'b001;
  assign for_1_for_for_k_2_0_1_sva_2 = nl_for_1_for_for_k_2_0_1_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_8_sva_2 = for_1_for_for_k_2_0_8_sva + 3'b001;
  assign for_1_for_for_k_2_0_8_sva_2 = nl_for_1_for_for_k_2_0_8_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_24_sva_2 = for_1_for_for_k_2_0_24_sva + 3'b001;
  assign for_1_for_for_k_2_0_24_sva_2 = nl_for_1_for_for_k_2_0_24_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_20_sva_2 = for_1_for_for_k_2_0_20_sva + 3'b001;
  assign for_1_for_for_k_2_0_20_sva_2 = nl_for_1_for_for_k_2_0_20_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_16_sva_2 = for_1_for_for_k_2_0_16_sva + 3'b001;
  assign for_1_for_for_k_2_0_16_sva_2 = nl_for_1_for_for_k_2_0_16_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_12_sva_2 = for_1_for_for_k_2_0_12_sva + 3'b001;
  assign for_1_for_for_k_2_0_12_sva_2 = nl_for_1_for_for_k_2_0_12_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_7_sva_2 = for_1_for_for_k_2_0_7_sva + 3'b001;
  assign for_1_for_for_k_2_0_7_sva_2 = nl_for_1_for_for_k_2_0_7_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_23_sva_2 = for_1_for_for_k_2_0_23_sva + 3'b001;
  assign for_1_for_for_k_2_0_23_sva_2 = nl_for_1_for_for_k_2_0_23_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_19_sva_2 = for_1_for_for_k_2_0_19_sva + 3'b001;
  assign for_1_for_for_k_2_0_19_sva_2 = nl_for_1_for_for_k_2_0_19_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_15_sva_2 = for_1_for_for_k_2_0_15_sva + 3'b001;
  assign for_1_for_for_k_2_0_15_sva_2 = nl_for_1_for_for_k_2_0_15_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_11_sva_2 = for_1_for_for_k_2_0_11_sva + 3'b001;
  assign for_1_for_for_k_2_0_11_sva_2 = nl_for_1_for_for_k_2_0_11_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_6_sva_2 = for_1_for_for_k_2_0_6_sva + 3'b001;
  assign for_1_for_for_k_2_0_6_sva_2 = nl_for_1_for_for_k_2_0_6_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_22_sva_2 = for_1_for_for_k_2_0_22_sva + 3'b001;
  assign for_1_for_for_k_2_0_22_sva_2 = nl_for_1_for_for_k_2_0_22_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_18_sva_2 = for_1_for_for_k_2_0_18_sva + 3'b001;
  assign for_1_for_for_k_2_0_18_sva_2 = nl_for_1_for_for_k_2_0_18_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_14_sva_2 = for_1_for_for_k_2_0_14_sva + 3'b001;
  assign for_1_for_for_k_2_0_14_sva_2 = nl_for_1_for_for_k_2_0_14_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_10_sva_2 = for_1_for_for_k_2_0_10_sva + 3'b001;
  assign for_1_for_for_k_2_0_10_sva_2 = nl_for_1_for_for_k_2_0_10_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_5_sva_2 = for_1_for_for_k_2_0_5_sva + 3'b001;
  assign for_1_for_for_k_2_0_5_sva_2 = nl_for_1_for_for_k_2_0_5_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_21_sva_2 = for_1_for_for_k_2_0_21_sva + 3'b001;
  assign for_1_for_for_k_2_0_21_sva_2 = nl_for_1_for_for_k_2_0_21_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_17_sva_2 = for_1_for_for_k_2_0_17_sva + 3'b001;
  assign for_1_for_for_k_2_0_17_sva_2 = nl_for_1_for_for_k_2_0_17_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_13_sva_2 = for_1_for_for_k_2_0_13_sva + 3'b001;
  assign for_1_for_for_k_2_0_13_sva_2 = nl_for_1_for_for_k_2_0_13_sva_2[2:0];
  assign nl_for_1_for_for_k_2_0_9_sva_2 = for_1_for_for_k_2_0_9_sva + 3'b001;
  assign for_1_for_for_k_2_0_9_sva_2 = nl_for_1_for_for_k_2_0_9_sva_2[2:0];
  assign for_1_5_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1 = MUX_v_16_8_2x1x2x3((a_value_value_sva[399:384]),
      (a_value_value_sva[335:320]), (a_value_value_sva[351:336]), (a_value_value_sva[367:352]),
      (a_value_value_sva[383:368]), {(~ (for_1_for_for_k_2_0_1_sva[2])) , (for_1_for_for_k_2_0_1_sva[1:0])});
  assign nl_for_1_1_for_for_acc_7_nl = for_1_for_for_k_2_0_5_sva + conv_u2u_1_3(for_1_for_for_k_2_0_5_sva[2])
      + 3'b001;
  assign for_1_1_for_for_acc_7_nl = nl_for_1_1_for_for_acc_7_nl[2:0];
  assign for_1_1_for_5_for_slc_b_value_value_16_15_0_ncse_sva_1 = MUX_v_16_25_2x0x1x2x3((b_value_value_sva[79:64]),
      (b_value_value_sva[95:80]), (b_value_value_sva[111:96]), (b_value_value_sva[127:112]),
      (b_value_value_sva[143:128]), (b_value_value_sva[159:144]), (b_value_value_sva[175:160]),
      (b_value_value_sva[191:176]), (b_value_value_sva[207:192]), (b_value_value_sva[223:208]),
      (b_value_value_sva[239:224]), (b_value_value_sva[255:240]), (b_value_value_sva[271:256]),
      (b_value_value_sva[287:272]), (b_value_value_sva[303:288]), (b_value_value_sva[319:304]),
      (b_value_value_sva[335:320]), (b_value_value_sva[351:336]), (b_value_value_sva[367:352]),
      (b_value_value_sva[383:368]), (b_value_value_sva[399:384]), {(for_1_1_for_for_acc_7_nl)
      , (for_1_for_for_k_2_0_5_sva[1:0])});
  assign nl_for_1_for_for_acc_19_nl = conv_u2u_1_3(for_1_for_for_acc_18_psp_1[2])
      + for_1_for_for_k_2_0_21_sva;
  assign for_1_for_for_acc_19_nl = nl_for_1_for_for_acc_19_nl[2:0];
  assign for_1_1_for_4_for_slc_b_value_value_16_15_0_ncse_sva_1 = MUX_v_16_24_2x0x1x2((b_value_value_sva[63:48]),
      (b_value_value_sva[79:64]), (b_value_value_sva[95:80]), (b_value_value_sva[111:96]),
      (b_value_value_sva[127:112]), (b_value_value_sva[143:128]), (b_value_value_sva[159:144]),
      (b_value_value_sva[175:160]), (b_value_value_sva[191:176]), (b_value_value_sva[207:192]),
      (b_value_value_sva[223:208]), (b_value_value_sva[239:224]), (b_value_value_sva[255:240]),
      (b_value_value_sva[271:256]), (b_value_value_sva[287:272]), (b_value_value_sva[303:288]),
      (b_value_value_sva[319:304]), (b_value_value_sva[335:320]), (b_value_value_sva[351:336]),
      (b_value_value_sva[367:352]), (b_value_value_sva[383:368]), {(for_1_for_for_acc_19_nl)
      , (for_1_for_for_acc_18_psp_1[1:0])});
  assign nl_for_1_1_for_for_acc_nl = ({for_1_for_for_k_2_0_17_sva , 1'b0}) + conv_u2u_2_4(for_1_for_for_k_2_0_17_sva[2:1])
      + 4'b0001;
  assign for_1_1_for_for_acc_nl = nl_for_1_1_for_for_acc_nl[3:0];
  assign for_1_1_for_3_for_slc_b_value_value_16_15_0_ncse_sva_1 = MUX_v_16_24_2x0x1((b_value_value_sva[47:32]),
      (b_value_value_sva[63:48]), (b_value_value_sva[79:64]), (b_value_value_sva[95:80]),
      (b_value_value_sva[111:96]), (b_value_value_sva[127:112]), (b_value_value_sva[143:128]),
      (b_value_value_sva[159:144]), (b_value_value_sva[175:160]), (b_value_value_sva[191:176]),
      (b_value_value_sva[207:192]), (b_value_value_sva[223:208]), (b_value_value_sva[239:224]),
      (b_value_value_sva[255:240]), (b_value_value_sva[271:256]), (b_value_value_sva[287:272]),
      (b_value_value_sva[303:288]), (b_value_value_sva[319:304]), (b_value_value_sva[335:320]),
      (b_value_value_sva[351:336]), (b_value_value_sva[367:352]), (b_value_value_sva[383:368]),
      {(for_1_1_for_for_acc_nl) , (for_1_for_for_k_2_0_17_sva[0])});
  assign nl_for_1_1_for_2_for_acc_6_nl = ({for_1_for_for_k_2_0_13_sva , 2'b00}) +
      conv_u2u_3_5(for_1_for_for_k_2_0_13_sva) + 5'b00001;
  assign for_1_1_for_2_for_acc_6_nl = nl_for_1_1_for_2_for_acc_6_nl[4:0];
  assign for_1_1_for_2_for_slc_b_value_value_16_15_0_ncse_sva_1 = MUX_v_16_22_2x0((b_value_value_sva[31:16]),
      (b_value_value_sva[47:32]), (b_value_value_sva[63:48]), (b_value_value_sva[79:64]),
      (b_value_value_sva[95:80]), (b_value_value_sva[111:96]), (b_value_value_sva[127:112]),
      (b_value_value_sva[143:128]), (b_value_value_sva[159:144]), (b_value_value_sva[175:160]),
      (b_value_value_sva[191:176]), (b_value_value_sva[207:192]), (b_value_value_sva[223:208]),
      (b_value_value_sva[239:224]), (b_value_value_sva[255:240]), (b_value_value_sva[271:256]),
      (b_value_value_sva[287:272]), (b_value_value_sva[303:288]), (b_value_value_sva[319:304]),
      (b_value_value_sva[335:320]), (b_value_value_sva[351:336]), for_1_1_for_2_for_acc_6_nl);
  assign nl_for_1_1_for_for_acc_8_nl = conv_u2u_1_3(for_1_for_for_k_2_0_9_sva[2])
      + for_1_for_for_k_2_0_9_sva;
  assign for_1_1_for_for_acc_8_nl = nl_for_1_1_for_for_acc_8_nl[2:0];
  assign for_1_1_for_1_for_slc_b_value_value_16_15_0_ncse_sva_1 = MUX_v_16_24_2((b_value_value_sva[15:0]),
      (b_value_value_sva[31:16]), (b_value_value_sva[47:32]), (b_value_value_sva[63:48]),
      (b_value_value_sva[79:64]), (b_value_value_sva[95:80]), (b_value_value_sva[111:96]),
      (b_value_value_sva[127:112]), (b_value_value_sva[143:128]), (b_value_value_sva[159:144]),
      (b_value_value_sva[175:160]), (b_value_value_sva[191:176]), (b_value_value_sva[207:192]),
      (b_value_value_sva[223:208]), (b_value_value_sva[239:224]), (b_value_value_sva[255:240]),
      (b_value_value_sva[271:256]), (b_value_value_sva[287:272]), (b_value_value_sva[303:288]),
      (b_value_value_sva[319:304]), (b_value_value_sva[335:320]), (b_value_value_sva[351:336]),
      (b_value_value_sva[367:352]), (b_value_value_sva[383:368]), {(for_1_1_for_for_acc_8_nl)
      , (for_1_for_for_k_2_0_9_sva[1:0])});
  assign nl_for_1_4_for_1_for_acc_5_nl = for_1_for_for_k_2_0_12_sva + 3'b111;
  assign for_1_4_for_1_for_acc_5_nl = nl_for_1_4_for_1_for_acc_5_nl[2:0];
  assign for_1_4_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1 = MUX_v_16_8_2x4x5x6((a_value_value_sva[271:256]),
      (a_value_value_sva[287:272]), (a_value_value_sva[303:288]), (a_value_value_sva[319:304]),
      (a_value_value_sva[255:240]), for_1_4_for_1_for_acc_5_nl);
  assign nl_for_1_for_for_acc_nl = (for_1_for_for_k_2_0_11_sva[2:1]) + 2'b01;
  assign for_1_for_for_acc_nl = nl_for_1_for_for_acc_nl[1:0];
  assign for_1_3_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1 = MUX_v_16_8_2x0x1((a_value_value_sva[175:160]),
      (a_value_value_sva[191:176]), (a_value_value_sva[207:192]), (a_value_value_sva[223:208]),
      (a_value_value_sva[239:224]), (a_value_value_sva[255:240]), {(for_1_for_for_acc_nl)
      , (for_1_for_for_k_2_0_11_sva[0])});
  assign nl_for_1_2_for_1_for_acc_5_nl = for_1_for_for_k_2_0_10_sva + 3'b101;
  assign for_1_2_for_1_for_acc_5_nl = nl_for_1_2_for_1_for_acc_5_nl[2:0];
  assign for_1_2_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1 = MUX_v_16_8_2x2x3x4((a_value_value_sva[143:128]),
      (a_value_value_sva[159:144]), (a_value_value_sva[95:80]), (a_value_value_sva[111:96]),
      (a_value_value_sva[127:112]), for_1_2_for_1_for_acc_5_nl);
  assign for_1_1_for_1_for_slc_a_value_value_16_15_0_ncse_sva_1 = MUX_v_16_5_2((a_value_value_sva[15:0]),
      (a_value_value_sva[31:16]), (a_value_value_sva[47:32]), (a_value_value_sva[63:48]),
      (a_value_value_sva[79:64]), for_1_for_for_k_2_0_9_sva);
  assign nl_for_1_for_for_acc_18_psp_1 = for_1_for_for_k_2_0_21_sva + 3'b011;
  assign for_1_for_for_acc_18_psp_1 = nl_for_1_for_for_acc_18_psp_1[2:0];
  assign nl_for_1_1_for_1_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_9_sva_2)
      + 4'b1011;
  assign for_1_1_for_1_for_acc_nl = nl_for_1_1_for_1_for_acc_nl[3:0];
  assign nl_for_1_1_for_2_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_13_sva_2)
      + 4'b1011;
  assign for_1_1_for_2_for_acc_nl = nl_for_1_1_for_2_for_acc_nl[3:0];
  assign nl_for_1_1_for_3_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_17_sva_2)
      + 4'b1011;
  assign for_1_1_for_3_for_acc_nl = nl_for_1_1_for_3_for_acc_nl[3:0];
  assign nl_for_1_1_for_4_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_21_sva_2)
      + 4'b1011;
  assign for_1_1_for_4_for_acc_nl = nl_for_1_1_for_4_for_acc_nl[3:0];
  assign nl_for_1_1_for_5_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_5_sva_2)
      + 4'b1011;
  assign for_1_1_for_5_for_acc_nl = nl_for_1_1_for_5_for_acc_nl[3:0];
  assign nl_for_1_2_for_1_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_10_sva_2)
      + 4'b1011;
  assign for_1_2_for_1_for_acc_nl = nl_for_1_2_for_1_for_acc_nl[3:0];
  assign nl_for_1_2_for_2_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_14_sva_2)
      + 4'b1011;
  assign for_1_2_for_2_for_acc_nl = nl_for_1_2_for_2_for_acc_nl[3:0];
  assign nl_for_1_2_for_3_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_18_sva_2)
      + 4'b1011;
  assign for_1_2_for_3_for_acc_nl = nl_for_1_2_for_3_for_acc_nl[3:0];
  assign nl_for_1_2_for_4_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_22_sva_2)
      + 4'b1011;
  assign for_1_2_for_4_for_acc_nl = nl_for_1_2_for_4_for_acc_nl[3:0];
  assign nl_for_1_2_for_5_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_6_sva_2)
      + 4'b1011;
  assign for_1_2_for_5_for_acc_nl = nl_for_1_2_for_5_for_acc_nl[3:0];
  assign nl_for_1_3_for_1_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_11_sva_2)
      + 4'b1011;
  assign for_1_3_for_1_for_acc_nl = nl_for_1_3_for_1_for_acc_nl[3:0];
  assign nl_for_1_3_for_2_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_15_sva_2)
      + 4'b1011;
  assign for_1_3_for_2_for_acc_nl = nl_for_1_3_for_2_for_acc_nl[3:0];
  assign nl_for_1_3_for_3_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_19_sva_2)
      + 4'b1011;
  assign for_1_3_for_3_for_acc_nl = nl_for_1_3_for_3_for_acc_nl[3:0];
  assign nl_for_1_3_for_4_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_23_sva_2)
      + 4'b1011;
  assign for_1_3_for_4_for_acc_nl = nl_for_1_3_for_4_for_acc_nl[3:0];
  assign nl_for_1_3_for_5_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_7_sva_2)
      + 4'b1011;
  assign for_1_3_for_5_for_acc_nl = nl_for_1_3_for_5_for_acc_nl[3:0];
  assign nl_for_1_4_for_1_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_12_sva_2)
      + 4'b1011;
  assign for_1_4_for_1_for_acc_nl = nl_for_1_4_for_1_for_acc_nl[3:0];
  assign nl_for_1_4_for_2_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_16_sva_2)
      + 4'b1011;
  assign for_1_4_for_2_for_acc_nl = nl_for_1_4_for_2_for_acc_nl[3:0];
  assign nl_for_1_4_for_3_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_20_sva_2)
      + 4'b1011;
  assign for_1_4_for_3_for_acc_nl = nl_for_1_4_for_3_for_acc_nl[3:0];
  assign nl_for_1_4_for_4_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_24_sva_2)
      + 4'b1011;
  assign for_1_4_for_4_for_acc_nl = nl_for_1_4_for_4_for_acc_nl[3:0];
  assign nl_for_1_4_for_5_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_8_sva_2)
      + 4'b1011;
  assign for_1_4_for_5_for_acc_nl = nl_for_1_4_for_5_for_acc_nl[3:0];
  assign nl_for_1_5_for_1_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_1_sva_2)
      + 4'b1011;
  assign for_1_5_for_1_for_acc_nl = nl_for_1_5_for_1_for_acc_nl[3:0];
  assign nl_for_1_5_for_2_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_2_sva_2)
      + 4'b1011;
  assign for_1_5_for_2_for_acc_nl = nl_for_1_5_for_2_for_acc_nl[3:0];
  assign nl_for_1_5_for_3_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_3_sva_2)
      + 4'b1011;
  assign for_1_5_for_3_for_acc_nl = nl_for_1_5_for_3_for_acc_nl[3:0];
  assign nl_for_1_5_for_4_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_4_sva_2)
      + 4'b1011;
  assign for_1_5_for_4_for_acc_nl = nl_for_1_5_for_4_for_acc_nl[3:0];
  assign nl_for_1_5_for_5_for_acc_nl = conv_u2s_3_4(for_1_for_for_k_2_0_sva_2) +
      4'b1011;
  assign for_1_5_for_5_for_acc_nl = nl_for_1_5_for_5_for_acc_nl[3:0];
  assign for_1_for_for_and_21_tmp = (~((readslicef_4_1_3((for_1_1_for_1_for_acc_nl)))
      | (readslicef_4_1_3((for_1_1_for_2_for_acc_nl))))) & (~((readslicef_4_1_3((for_1_1_for_3_for_acc_nl)))
      | (readslicef_4_1_3((for_1_1_for_4_for_acc_nl))))) & (~((readslicef_4_1_3((for_1_1_for_5_for_acc_nl)))
      | (readslicef_4_1_3((for_1_2_for_1_for_acc_nl))))) & (~((readslicef_4_1_3((for_1_2_for_2_for_acc_nl)))
      | (readslicef_4_1_3((for_1_2_for_3_for_acc_nl))))) & (~((readslicef_4_1_3((for_1_2_for_4_for_acc_nl)))
      | (readslicef_4_1_3((for_1_2_for_5_for_acc_nl))))) & (~((readslicef_4_1_3((for_1_3_for_1_for_acc_nl)))
      | (readslicef_4_1_3((for_1_3_for_2_for_acc_nl))))) & (~((readslicef_4_1_3((for_1_3_for_3_for_acc_nl)))
      | (readslicef_4_1_3((for_1_3_for_4_for_acc_nl))))) & (~((readslicef_4_1_3((for_1_3_for_5_for_acc_nl)))
      | (readslicef_4_1_3((for_1_4_for_1_for_acc_nl))))) & (~((readslicef_4_1_3((for_1_4_for_2_for_acc_nl)))
      | (readslicef_4_1_3((for_1_4_for_3_for_acc_nl))) | (readslicef_4_1_3((for_1_4_for_4_for_acc_nl)))
      | (readslicef_4_1_3((for_1_4_for_5_for_acc_nl))) | (readslicef_4_1_3((for_1_5_for_1_for_acc_nl)))
      | (readslicef_4_1_3((for_1_5_for_2_for_acc_nl))) | (readslicef_4_1_3((for_1_5_for_3_for_acc_nl)))
      | (readslicef_4_1_3((for_1_5_for_4_for_acc_nl))) | (readslicef_4_1_3((for_1_5_for_5_for_acc_nl)))));
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      c_chan_rsci_idat_15_0 <= 16'b0000000000000000;
      c_chan_rsci_idat_31_16 <= 16'b0000000000000000;
      c_chan_rsci_idat_47_32 <= 16'b0000000000000000;
      c_chan_rsci_idat_63_48 <= 16'b0000000000000000;
      c_chan_rsci_idat_79_64 <= 16'b0000000000000000;
      c_chan_rsci_idat_95_80 <= 16'b0000000000000000;
      c_chan_rsci_idat_111_96 <= 16'b0000000000000000;
      c_chan_rsci_idat_127_112 <= 16'b0000000000000000;
      c_chan_rsci_idat_143_128 <= 16'b0000000000000000;
      c_chan_rsci_idat_159_144 <= 16'b0000000000000000;
      c_chan_rsci_idat_175_160 <= 16'b0000000000000000;
      c_chan_rsci_idat_191_176 <= 16'b0000000000000000;
      c_chan_rsci_idat_207_192 <= 16'b0000000000000000;
      c_chan_rsci_idat_223_208 <= 16'b0000000000000000;
      c_chan_rsci_idat_239_224 <= 16'b0000000000000000;
      c_chan_rsci_idat_255_240 <= 16'b0000000000000000;
      c_chan_rsci_idat_271_256 <= 16'b0000000000000000;
      c_chan_rsci_idat_287_272 <= 16'b0000000000000000;
      c_chan_rsci_idat_303_288 <= 16'b0000000000000000;
      c_chan_rsci_idat_319_304 <= 16'b0000000000000000;
      c_chan_rsci_idat_335_320 <= 16'b0000000000000000;
      c_chan_rsci_idat_351_336 <= 16'b0000000000000000;
      c_chan_rsci_idat_367_352 <= 16'b0000000000000000;
      c_chan_rsci_idat_383_368 <= 16'b0000000000000000;
      c_chan_rsci_idat_399_384 <= 16'b0000000000000000;
    end
    else if ( c_chan_and_cse ) begin
      c_chan_rsci_idat_15_0 <= for_1_for_tmp_9_sva_1_mx0w0;
      c_chan_rsci_idat_31_16 <= for_1_for_tmp_13_sva_1_mx0w0;
      c_chan_rsci_idat_47_32 <= for_1_for_tmp_17_sva_1_mx0w0;
      c_chan_rsci_idat_63_48 <= for_1_for_tmp_21_sva_1_mx0w0;
      c_chan_rsci_idat_79_64 <= for_1_for_tmp_5_sva_1_mx0w0;
      c_chan_rsci_idat_95_80 <= for_1_for_tmp_10_sva_1_mx0w0;
      c_chan_rsci_idat_111_96 <= for_1_for_tmp_14_sva_1_mx0w0;
      c_chan_rsci_idat_127_112 <= for_1_for_tmp_18_sva_1_mx0w0;
      c_chan_rsci_idat_143_128 <= for_1_for_tmp_22_sva_1_mx0w0;
      c_chan_rsci_idat_159_144 <= for_1_for_tmp_6_sva_1_mx0w0;
      c_chan_rsci_idat_175_160 <= for_1_for_tmp_11_sva_1_mx0w0;
      c_chan_rsci_idat_191_176 <= for_1_for_tmp_15_sva_1_mx0w0;
      c_chan_rsci_idat_207_192 <= for_1_for_tmp_19_sva_1_mx0w0;
      c_chan_rsci_idat_223_208 <= for_1_for_tmp_23_sva_1_mx0w0;
      c_chan_rsci_idat_239_224 <= for_1_for_tmp_7_sva_1_mx0w0;
      c_chan_rsci_idat_255_240 <= for_1_for_tmp_12_sva_1_mx0w0;
      c_chan_rsci_idat_271_256 <= for_1_for_tmp_16_sva_1_mx0w0;
      c_chan_rsci_idat_287_272 <= for_1_for_tmp_20_sva_1_mx0w0;
      c_chan_rsci_idat_303_288 <= for_1_for_tmp_24_sva_1_mx0w0;
      c_chan_rsci_idat_319_304 <= for_1_for_tmp_8_sva_1_mx0w0;
      c_chan_rsci_idat_335_320 <= for_1_for_tmp_1_sva_1_mx0w0;
      c_chan_rsci_idat_351_336 <= for_1_for_tmp_2_sva_1_mx0w0;
      c_chan_rsci_idat_367_352 <= for_1_for_tmp_3_sva_1_mx0w0;
      c_chan_rsci_idat_383_368 <= for_1_for_tmp_4_sva_1_mx0w0;
      c_chan_rsci_idat_399_384 <= for_1_for_tmp_sva_1_mx0w0;
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      reg_c_chan_rsci_ivld_run_psct_cse <= 1'b0;
      reg_b_chan_rsci_irdy_run_psct_cse <= 1'b0;
      for_1_for_for_k_2_0_sva <= 3'b000;
      for_1_for_tmp_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_4_sva <= 3'b000;
      for_1_for_tmp_4_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_3_sva <= 3'b000;
      for_1_for_tmp_3_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_2_sva <= 3'b000;
      for_1_for_tmp_2_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_1_sva <= 3'b000;
      for_1_for_tmp_1_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_8_sva <= 3'b000;
      for_1_for_tmp_8_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_24_sva <= 3'b000;
      for_1_for_tmp_24_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_20_sva <= 3'b000;
      for_1_for_tmp_20_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_16_sva <= 3'b000;
      for_1_for_tmp_16_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_12_sva <= 3'b000;
      for_1_for_tmp_12_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_7_sva <= 3'b000;
      for_1_for_tmp_7_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_23_sva <= 3'b000;
      for_1_for_tmp_23_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_19_sva <= 3'b000;
      for_1_for_tmp_19_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_15_sva <= 3'b000;
      for_1_for_tmp_15_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_11_sva <= 3'b000;
      for_1_for_tmp_11_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_6_sva <= 3'b000;
      for_1_for_tmp_6_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_22_sva <= 3'b000;
      for_1_for_tmp_22_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_18_sva <= 3'b000;
      for_1_for_tmp_18_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_14_sva <= 3'b000;
      for_1_for_tmp_14_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_10_sva <= 3'b000;
      for_1_for_tmp_10_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_5_sva <= 3'b000;
      for_1_for_tmp_5_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_21_sva <= 3'b000;
      for_1_for_tmp_21_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_17_sva <= 3'b000;
      for_1_for_tmp_17_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_13_sva <= 3'b000;
      for_1_for_tmp_13_sva <= 16'b0000000000000000;
      for_1_for_for_k_2_0_9_sva <= 3'b000;
      for_1_for_tmp_9_sva <= 16'b0000000000000000;
    end
    else if ( run_wen ) begin
      reg_c_chan_rsci_ivld_run_psct_cse <= for_1_for_for_and_21_tmp & (fsm_output[2]);
      reg_b_chan_rsci_irdy_run_psct_cse <= ~((fsm_output[2:1]!=2'b00));
      for_1_for_for_k_2_0_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_sva_2, (fsm_output[2]));
      for_1_for_tmp_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_4_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_4_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_4_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_4_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_3_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_3_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_3_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_3_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_2_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_2_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_2_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_2_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_1_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_1_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_1_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_1_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_8_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_8_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_8_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_8_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_24_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_24_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_24_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_24_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_20_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_20_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_20_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_20_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_16_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_16_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_16_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_16_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_12_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_12_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_12_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_12_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_7_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_7_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_7_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_7_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_23_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_23_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_23_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_23_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_19_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_19_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_19_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_19_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_15_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_15_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_15_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_15_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_11_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_11_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_11_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_11_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_6_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_6_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_6_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_6_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_22_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_22_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_22_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_22_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_18_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_18_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_18_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_18_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_14_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_14_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_14_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_14_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_10_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_10_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_10_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_10_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_5_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_5_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_5_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_5_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_21_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_21_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_21_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_21_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_17_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_17_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_17_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_17_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_13_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_13_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_13_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_13_sva_1_mx0w0,
          (fsm_output[2]));
      for_1_for_for_k_2_0_9_sva <= MUX_v_3_2_2(3'b000, for_1_for_for_k_2_0_9_sva_2,
          (fsm_output[2]));
      for_1_for_tmp_9_sva <= MUX_v_16_2_2(16'b0000000000000000, for_1_for_tmp_9_sva_1_mx0w0,
          (fsm_output[2]));
    end
  end
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      a_value_value_sva <= 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
      b_value_value_sva <= 400'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( a_value_value_and_cse ) begin
      a_value_value_sva <= a_chan_rsci_idat_mxwt;
      b_value_value_sva <= b_chan_rsci_idat_mxwt;
    end
  end

  function automatic [15:0] MUX_v_16_22_2x0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [4:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      default : begin
        result = input_21;
      end
    endcase
    MUX_v_16_22_2x0 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_24_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [4:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      5'b00000 : begin
        result = input_0;
      end
      5'b00001 : begin
        result = input_1;
      end
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      default : begin
        result = input_23;
      end
    endcase
    MUX_v_16_24_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_24_2x0x1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [4:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      5'b00010 : begin
        result = input_2;
      end
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      default : begin
        result = input_23;
      end
    endcase
    MUX_v_16_24_2x0x1 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_24_2x0x1x2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [4:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      5'b00011 : begin
        result = input_3;
      end
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      default : begin
        result = input_23;
      end
    endcase
    MUX_v_16_24_2x0x1x2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_25_2x0x1x2x3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [15:0] input_8;
    input [15:0] input_9;
    input [15:0] input_10;
    input [15:0] input_11;
    input [15:0] input_12;
    input [15:0] input_13;
    input [15:0] input_14;
    input [15:0] input_15;
    input [15:0] input_16;
    input [15:0] input_17;
    input [15:0] input_18;
    input [15:0] input_19;
    input [15:0] input_20;
    input [15:0] input_21;
    input [15:0] input_22;
    input [15:0] input_23;
    input [15:0] input_24;
    input [4:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      5'b00100 : begin
        result = input_4;
      end
      5'b00101 : begin
        result = input_5;
      end
      5'b00110 : begin
        result = input_6;
      end
      5'b00111 : begin
        result = input_7;
      end
      5'b01000 : begin
        result = input_8;
      end
      5'b01001 : begin
        result = input_9;
      end
      5'b01010 : begin
        result = input_10;
      end
      5'b01011 : begin
        result = input_11;
      end
      5'b01100 : begin
        result = input_12;
      end
      5'b01101 : begin
        result = input_13;
      end
      5'b01110 : begin
        result = input_14;
      end
      5'b01111 : begin
        result = input_15;
      end
      5'b10000 : begin
        result = input_16;
      end
      5'b10001 : begin
        result = input_17;
      end
      5'b10010 : begin
        result = input_18;
      end
      5'b10011 : begin
        result = input_19;
      end
      5'b10100 : begin
        result = input_20;
      end
      5'b10101 : begin
        result = input_21;
      end
      5'b10110 : begin
        result = input_22;
      end
      5'b10111 : begin
        result = input_23;
      end
      default : begin
        result = input_24;
      end
    endcase
    MUX_v_16_25_2x0x1x2x3 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_2_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [0:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_16_2_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_5_2;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [2:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      default : begin
        result = input_4;
      end
    endcase
    MUX_v_16_5_2 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_8_2x0x1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [2:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_16_8_2x0x1 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_8_2x1x2x3;
    input [15:0] input_0;
    input [15:0] input_4;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [2:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_16_8_2x1x2x3 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_8_2x2x3x4;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_5;
    input [15:0] input_6;
    input [15:0] input_7;
    input [2:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_16_8_2x2x3x4 = result;
  end
  endfunction


  function automatic [15:0] MUX_v_16_8_2x4x5x6;
    input [15:0] input_0;
    input [15:0] input_1;
    input [15:0] input_2;
    input [15:0] input_3;
    input [15:0] input_7;
    input [2:0] sel;
    reg [15:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_16_8_2x4x5x6 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_4_1_3;
    input [3:0] vector;
    reg [3:0] tmp;
  begin
    tmp = vector >> 3;
    readslicef_4_1_3 = tmp[0:0];
  end
  endfunction


  function automatic [3:0] conv_u2s_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2s_3_4 =  {1'b0, vector};
  end
  endfunction


  function automatic [2:0] conv_u2u_1_3 ;
    input [0:0]  vector ;
  begin
    conv_u2u_1_3 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_2_4 ;
    input [1:0]  vector ;
  begin
    conv_u2u_2_4 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [4:0] conv_u2u_3_5 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_5 = {{2{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult_struct
// ------------------------------------------------------------------


module MatMult_struct (
  clk, arst_n, a_chan_rsc_dat_value, a_chan_rsc_vld, a_chan_rsc_rdy, b_chan_rsc_dat_value,
      b_chan_rsc_vld, b_chan_rsc_rdy, c_chan_rsc_dat_value, c_chan_rsc_vld, c_chan_rsc_rdy
);
  input clk;
  input arst_n;
  input [399:0] a_chan_rsc_dat_value;
  input a_chan_rsc_vld;
  output a_chan_rsc_rdy;
  input [399:0] b_chan_rsc_dat_value;
  input b_chan_rsc_vld;
  output b_chan_rsc_rdy;
  output [399:0] c_chan_rsc_dat_value;
  output c_chan_rsc_vld;
  input c_chan_rsc_rdy;


  // Interconnect Declarations
  wire [399:0] c_chan_rsc_dat;


  // Interconnect Declarations for Component Instantiations 
  MatMult_run MatMult_run_inst (
      .clk(clk),
      .arst_n(arst_n),
      .a_chan_rsc_dat(a_chan_rsc_dat_value),
      .a_chan_rsc_vld(a_chan_rsc_vld),
      .a_chan_rsc_rdy(a_chan_rsc_rdy),
      .b_chan_rsc_dat(b_chan_rsc_dat_value),
      .b_chan_rsc_vld(b_chan_rsc_vld),
      .b_chan_rsc_rdy(b_chan_rsc_rdy),
      .c_chan_rsc_dat(c_chan_rsc_dat),
      .c_chan_rsc_vld(c_chan_rsc_vld),
      .c_chan_rsc_rdy(c_chan_rsc_rdy)
    );
  assign c_chan_rsc_dat_value = c_chan_rsc_dat;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    MatMult
// ------------------------------------------------------------------


module MatMult (
  clk, arst_n, a_chan_rsc_dat, a_chan_rsc_vld, a_chan_rsc_rdy, b_chan_rsc_dat, b_chan_rsc_vld,
      b_chan_rsc_rdy, c_chan_rsc_dat, c_chan_rsc_vld, c_chan_rsc_rdy
);
  input clk;
  input arst_n;
  input [399:0] a_chan_rsc_dat;
  input a_chan_rsc_vld;
  output a_chan_rsc_rdy;
  input [399:0] b_chan_rsc_dat;
  input b_chan_rsc_vld;
  output b_chan_rsc_rdy;
  output [399:0] c_chan_rsc_dat;
  output c_chan_rsc_vld;
  input c_chan_rsc_rdy;


  // Interconnect Declarations
  wire [399:0] c_chan_rsc_dat_value;


  // Interconnect Declarations for Component Instantiations 
  MatMult_struct MatMult_struct_inst (
      .clk(clk),
      .arst_n(arst_n),
      .a_chan_rsc_dat_value(a_chan_rsc_dat),
      .a_chan_rsc_vld(a_chan_rsc_vld),
      .a_chan_rsc_rdy(a_chan_rsc_rdy),
      .b_chan_rsc_dat_value(b_chan_rsc_dat),
      .b_chan_rsc_vld(b_chan_rsc_vld),
      .b_chan_rsc_rdy(b_chan_rsc_rdy),
      .c_chan_rsc_dat_value(c_chan_rsc_dat_value),
      .c_chan_rsc_vld(c_chan_rsc_vld),
      .c_chan_rsc_rdy(c_chan_rsc_rdy)
    );
  assign c_chan_rsc_dat = c_chan_rsc_dat_value;
endmodule



